module work1 (clk_in, clk_out, reset);
parameter n = 7;
input clk_in, reset;
output clk_out;

reg clk1, clk2;
reg [7:0] count;

always @(posedge clk_in or posedge reset) begin
	if (reset) begin
		count <= n-1;
	end
	else if (count == n-1)
		count <= 0;
	else
		count <= count + 1;
end

always @(posedge clk_in or posedge reset) begin
	if (reset) 
		clk1 <= 1;
	else if (count == n-1)
		clk1 <= ~clk1;
	else
		clk1 <= clk1;
end

always @(negedge clk_in or posedge reset) begin
	if (reset)
		clk2 <= 1;
	else if (count == (n-1)/2)
		clk2 <= ~clk2;
	else 
		clk2 <= clk2;
end

assign clk_out = clk1 ^ clk2;

endmodule
