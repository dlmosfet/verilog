library verilog;
use verilog.vl_types.all;
entity work1_vlg_vec_tst is
end work1_vlg_vec_tst;
